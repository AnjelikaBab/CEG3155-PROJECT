library verilog;
use verilog.vl_types.all;
entity baudRateGenerator_vlg_vec_tst is
end baudRateGenerator_vlg_vec_tst;
