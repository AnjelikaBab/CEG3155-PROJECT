library verilog;
use verilog.vl_types.all;
entity uartTopLevel_vlg_vec_tst is
end uartTopLevel_vlg_vec_tst;
